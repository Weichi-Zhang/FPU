`ifndef __PARAMS_VH__
`define __PARAMS_VH__

parameter EXPWIDTH = 8;
parameter SIGWIDTH = 24;
parameter XLEN = 32;

`endif
