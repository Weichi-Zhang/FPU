`ifndef __PARAMS_VH__
`define __PARAMS_VH__

parameter EXPWIDTH = 8;
parameter SIGWIDTH = 24;
parameter XLEN = 32;
parameter FLEN = 32;
parameter VIR_REG_ADDR_WIDTH = 6;

`endif
